module SignalGenerator(
    input wire clk
);

endmodule