module uart_tb(
    
);